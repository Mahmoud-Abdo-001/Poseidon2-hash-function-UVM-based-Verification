package crypto_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "crypto_seq_item.sv"   
    `include "crypto_config_obj.sv" 

    `include "sequencer.sv"
    `include "random_sequence.sv"

    `include "crypto_driver.sv"
    `include "crypto_monitor.sv"
    `include "crypto_agent.sv"
    `include "crypto_scoreboard.sv"
    `include "crypto_coverage_collector.sv"

    `include "crypto_environment.sv"
    `include "crypto_test.sv"

endpackage